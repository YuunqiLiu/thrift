

module top;


    bit                 var_bit         ;
    byte                var_byte        ;
    shortint            var_shortint    ;
    int                 var_int         ;
    longint             var_longint     ;
    byte unsigned       var_u_byte      ;
    shortint unsigned   var_u_shortint  ;
    int unsigned        var_u_int       ;
    longint unsigned    var_u_longint   ;
    real                var_real        ;
    shortreal           var_shortreal   ;
    string              var_string      ;

    initial begin

    end


endmodule